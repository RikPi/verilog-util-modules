module spi_master_cu #(
    parameter fifo_depth = 8
) (
    input wire clk,
    input wire aReset,
    input wire i_stream_in,
    output wire o_stream_out,
    input wire i_datapck_in,
    output wire o_datapck_out

);
    
endmodule